
`ifndef TEST_PACKAGE
`define TEST_PACKAGE
package symbol_gen_test_pkg;


 import uvm_pkg::*;
 `include "uvm_macros.svh"

 import global_defs_pkg::*;

 // TestBench specific imports

 import symbol_gen_reg_block_pkg::symbol_gen_reg_block;
 import symbol_gen_agent_pkg::*;
 import symbol_gen_agent_seq_pkg::*;
 import reset_agent_pkg::*;
 import reset_agent_seq_pkg::*;
 import clock_agent_pkg::*;
 import clock_agent_seq_pkg::*;
 import wb_agent_pkg::*;
 import wb_agent_seq_pkg::*;
 import symbol_gen_vseq_pkg::*;
 import symbol_gen_env_pkg::*;



 `include "symbol_gen_base_test.svh"
 `include "symbol_gen_base_test_user.svh"

 `include "symbol_gen_write_read_test.svh"




endpackage
`endif
