
`ifndef clock_agent_defines
`define clock_agent_defines

//Defines specific to this agent
`endif
