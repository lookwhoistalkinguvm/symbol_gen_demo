
`ifndef symbol_gen_agent_defines
`define symbol_gen_agent_defines

//Defines specific to this agent
`endif
