
`ifndef wb_agent_defines
`define wb_agent_defines

//Defines specific to this agent
`endif
