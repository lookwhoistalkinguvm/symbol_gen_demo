
`ifndef reset_agent_defines
`define reset_agent_defines

//Defines specific to this agent
`endif
