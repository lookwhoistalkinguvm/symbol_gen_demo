
`ifndef symbol_gen_vseq_pkg;
`define symbol_gen_vseq_pkg;

package symbol_gen_vseq_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import global_defs_pkg::*;


// Imports

 import symbol_gen_agent_pkg::*;
 import symbol_gen_agent_seq_pkg::*;
 import reset_agent_pkg::*;
 import reset_agent_seq_pkg::*;
 import clock_agent_pkg::*;
 import clock_agent_seq_pkg::*;
 import wb_agent_pkg::*;
 import wb_agent_seq_pkg::*;
 import symbol_gen_reg_block_pkg::symbol_gen_reg_block;
 import symbol_gen_env_pkg::*;


// Includes

 `include "symbol_gen_base_vseq.svh"
 `include "symbol_gen_base_user_vseq.svh"
 `include "symbol_gen_write_read_vseq.svh"


endpackage
`endif
