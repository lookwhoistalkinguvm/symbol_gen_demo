
`ifndef symbol_gen_env_config_user
`define symbol_gen_env_config_user

class symbol_gen_env_config_user extends symbol_gen_env_config;
`uvm_object_utils(symbol_gen_env_config_user)


endclass
`endif
