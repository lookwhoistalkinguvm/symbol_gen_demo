

package symbol_gen_reg_block_pkg;

 import uvm_pkg::*;
 `include "uvm_macros.svh"


 `include "PRERhi.svh"
 `include "TXR.svh"
 `include "RXR.svh"
 `include "CR.svh"
 `include "CTR.svh"
 `include "SR.svh"
 `include "PRERlo.svh"


 `include "symbol_gen_reg_block.svh"




endpackage
