
`ifndef symbol_gen_agent_seq_pkg;
`define symbol_gen_agent_seq_pkg;

package symbol_gen_agent_seq_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import global_defs_pkg::*;

 import symbol_gen_reg_block_pkg::symbol_gen_reg_block;
 import symbol_gen_agent_pkg::*;


// Symbol Sequences

 `include "symbol_gen_base_seq.svh"
 `include "symbol_gen_blocking_symbol_seq.svh"
 `include "symbol_gen_idle_symbol_seq.svh"
 `include "symbol_gen_slave_start_symbol_seq.svh"
 `include "symbol_gen_slave_listen_bit_symbol_seq.svh"
 `include "symbol_gen_slave_drive_bit_low_symbol_seq.svh"
 `include "monitor_symbol_gen_start_symbol_seq.svh"
 `include "monitor_symbol_gen_listen_bit_symbol_seq.svh"
 `include "monitor_symbol_gen_drive_bit_low_symbol_seq.svh"


// Sequences

 `include "symbol_gen_slave_address_seq.svh"




endpackage

`endif
